library verilog;
use verilog.vl_types.all;
entity ddr2_phy is
    port(
        pll_ref_clk     : in     vl_logic;
        global_reset_n  : in     vl_logic;
        soft_reset_n    : in     vl_logic;
        ctl_dqs_burst   : in     vl_logic_vector(1 downto 0);
        ctl_wdata_valid : in     vl_logic_vector(1 downto 0);
        ctl_wdata       : in     vl_logic_vector(31 downto 0);
        ctl_dm          : in     vl_logic_vector(3 downto 0);
        ctl_addr        : in     vl_logic_vector(12 downto 0);
        ctl_ba          : in     vl_logic_vector(2 downto 0);
        ctl_cas_n       : in     vl_logic_vector(0 downto 0);
        ctl_cke         : in     vl_logic_vector(0 downto 0);
        ctl_cs_n        : in     vl_logic_vector(0 downto 0);
        ctl_odt         : in     vl_logic_vector(0 downto 0);
        ctl_ras_n       : in     vl_logic_vector(0 downto 0);
        ctl_we_n        : in     vl_logic_vector(0 downto 0);
        ctl_rst_n       : in     vl_logic_vector(0 downto 0);
        ctl_mem_clk_disable: in     vl_logic_vector(0 downto 0);
        ctl_doing_rd    : in     vl_logic_vector(1 downto 0);
        ctl_cal_req     : in     vl_logic;
        ctl_cal_byte_lane_sel_n: in     vl_logic_vector(1 downto 0);
        dbg_clk         : in     vl_logic;
        dbg_reset_n     : in     vl_logic;
        dbg_addr        : in     vl_logic_vector(12 downto 0);
        dbg_wr          : in     vl_logic;
        dbg_rd          : in     vl_logic;
        dbg_cs          : in     vl_logic;
        dbg_wr_data     : in     vl_logic_vector(31 downto 0);
        reset_request_n : out    vl_logic;
        ctl_clk         : out    vl_logic;
        ctl_reset_n     : out    vl_logic;
        ctl_wlat        : out    vl_logic_vector(4 downto 0);
        ctl_rdata       : out    vl_logic_vector(31 downto 0);
        ctl_rdata_valid : out    vl_logic_vector(0 downto 0);
        ctl_rlat        : out    vl_logic_vector(4 downto 0);
        ctl_cal_success : out    vl_logic;
        ctl_cal_fail    : out    vl_logic;
        ctl_cal_warning : out    vl_logic;
        mem_addr        : out    vl_logic_vector(12 downto 0);
        mem_ba          : out    vl_logic_vector(2 downto 0);
        mem_cas_n       : out    vl_logic;
        mem_cke         : out    vl_logic_vector(0 downto 0);
        mem_cs_n        : out    vl_logic_vector(0 downto 0);
        mem_dm          : out    vl_logic_vector(1 downto 0);
        mem_odt         : out    vl_logic_vector(0 downto 0);
        mem_ras_n       : out    vl_logic;
        mem_we_n        : out    vl_logic;
        mem_reset_n     : out    vl_logic;
        dbg_rd_data     : out    vl_logic_vector(31 downto 0);
        dbg_waitrequest : out    vl_logic;
        aux_half_rate_clk: out    vl_logic;
        aux_full_rate_clk: out    vl_logic;
        mem_clk         : inout  vl_logic_vector(0 downto 0);
        mem_clk_n       : inout  vl_logic_vector(0 downto 0);
        mem_dq          : inout  vl_logic_vector(15 downto 0);
        mem_dqs         : inout  vl_logic_vector(1 downto 0);
        mem_dqs_n       : inout  vl_logic_vector(1 downto 0)
    );
end ddr2_phy;
