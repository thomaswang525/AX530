library verilog;
use verilog.vl_types.all;
entity ddr2_phy_alt_mem_phy_mux is
    generic(
        LOCAL_IF_AWIDTH : integer := 26;
        LOCAL_IF_DWIDTH : integer := 256;
        LOCAL_BURST_LEN_BITS: integer := 1;
        MEM_IF_DQ_PER_DQS: integer := 8;
        MEM_IF_DWIDTH   : integer := 64
    );
    port(
        phy_clk_1x      : in     vl_logic;
        reset_phy_clk_1x_n: in     vl_logic;
        ctl_address     : out    vl_logic_vector;
        ctl_read_req    : out    vl_logic;
        ctl_wdata       : out    vl_logic_vector;
        ctl_write_req   : out    vl_logic;
        ctl_size        : out    vl_logic_vector;
        ctl_be          : out    vl_logic_vector;
        ctl_refresh_req : out    vl_logic;
        ctl_burstbegin  : out    vl_logic;
        ctl_ready       : in     vl_logic;
        ctl_wdata_req   : in     vl_logic;
        ctl_rdata       : in     vl_logic_vector;
        ctl_rdata_valid : in     vl_logic;
        ctl_refresh_ack : in     vl_logic;
        ctl_init_done   : in     vl_logic;
        ctl_usr_mode_rdy: in     vl_logic;
        local_address   : in     vl_logic_vector;
        local_read_req  : in     vl_logic;
        local_wdata     : in     vl_logic_vector;
        local_write_req : in     vl_logic;
        local_size      : in     vl_logic_vector;
        local_be        : in     vl_logic_vector;
        local_refresh_req: in     vl_logic;
        local_burstbegin: in     vl_logic;
        mux_seq_controller_ready: out    vl_logic;
        mux_seq_wdata_req: out    vl_logic;
        seq_mux_address : in     vl_logic_vector;
        seq_mux_read_req: in     vl_logic;
        seq_mux_wdata   : in     vl_logic_vector;
        seq_mux_write_req: in     vl_logic;
        seq_mux_size    : in     vl_logic_vector;
        seq_mux_be      : in     vl_logic_vector;
        seq_mux_refresh_req: in     vl_logic;
        seq_mux_burstbegin: in     vl_logic;
        local_autopch_req: in     vl_logic;
        local_powerdn_req: in     vl_logic;
        local_self_rfsh_req: in     vl_logic;
        local_powerdn_ack: out    vl_logic;
        local_self_rfsh_ack: out    vl_logic;
        ctl_autopch_req : out    vl_logic;
        ctl_powerdn_req : out    vl_logic;
        ctl_self_rfsh_req: out    vl_logic;
        ctl_powerdn_ack : in     vl_logic;
        ctl_self_rfsh_ack: in     vl_logic;
        local_ready     : out    vl_logic;
        local_wdata_req : out    vl_logic;
        local_init_done : out    vl_logic;
        local_rdata     : out    vl_logic_vector;
        local_rdata_valid: out    vl_logic;
        local_refresh_ack: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOCAL_IF_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_IF_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_BURST_LEN_BITS : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQ_PER_DQS : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DWIDTH : constant is 1;
end ddr2_phy_alt_mem_phy_mux;
