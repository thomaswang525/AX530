library verilog;
use verilog.vl_types.all;
entity ddr2_phy_alt_mem_phy_seq_wrapper is
    port(
        phy_clk_1x      : in     vl_logic;
        reset_phy_clk_1x_n: in     vl_logic;
        ctl_cal_success : out    vl_logic;
        ctl_cal_fail    : out    vl_logic;
        ctl_cal_warning : out    vl_logic;
        ctl_cal_req     : in     vl_logic;
        int_RANK_HAS_ADDR_SWAP: in     vl_logic_vector(0 downto 0);
        ctl_cal_byte_lane_sel_n: in     vl_logic_vector(1 downto 0);
        seq_pll_inc_dec_n: out    vl_logic;
        seq_pll_start_reconfig: out    vl_logic;
        seq_pll_select  : out    vl_logic_vector(2 downto 0);
        phs_shft_busy   : in     vl_logic;
        pll_resync_clk_index: in     vl_logic_vector(2 downto 0);
        pll_measure_clk_index: in     vl_logic_vector(2 downto 0);
        sc_clk_dp       : out    vl_logic_vector(1 downto 0);
        scan_enable_dqs_config: out    vl_logic_vector(1 downto 0);
        scan_update     : out    vl_logic_vector(1 downto 0);
        scan_din        : out    vl_logic_vector(1 downto 0);
        scan_enable_ck  : out    vl_logic_vector(0 downto 0);
        scan_enable_dqs : out    vl_logic_vector(1 downto 0);
        scan_enable_dqsn: out    vl_logic_vector(1 downto 0);
        scan_enable_dq  : out    vl_logic_vector(15 downto 0);
        scan_enable_dm  : out    vl_logic_vector(1 downto 0);
        hr_rsc_clk      : in     vl_logic;
        seq_ac_addr     : out    vl_logic_vector(12 downto 0);
        seq_ac_ba       : out    vl_logic_vector(2 downto 0);
        seq_ac_cas_n    : out    vl_logic_vector(0 downto 0);
        seq_ac_ras_n    : out    vl_logic_vector(0 downto 0);
        seq_ac_we_n     : out    vl_logic_vector(0 downto 0);
        seq_ac_cke      : out    vl_logic_vector(0 downto 0);
        seq_ac_cs_n     : out    vl_logic_vector(0 downto 0);
        seq_ac_odt      : out    vl_logic_vector(0 downto 0);
        seq_ac_rst_n    : out    vl_logic_vector(0 downto 0);
        seq_ac_sel      : out    vl_logic;
        seq_mem_clk_disable: out    vl_logic;
        ctl_add_1t_ac_lat_internal: out    vl_logic;
        ctl_add_1t_odt_lat_internal: out    vl_logic;
        ctl_add_intermediate_regs_internal: out    vl_logic;
        seq_rdv_doing_rd: out    vl_logic_vector(1 downto 0);
        seq_rdp_reset_req_n: out    vl_logic;
        seq_rdp_inc_read_lat_1x: out    vl_logic_vector(1 downto 0);
        seq_rdp_dec_read_lat_1x: out    vl_logic_vector(1 downto 0);
        ctl_rdata       : in     vl_logic_vector(31 downto 0);
        int_rdata_valid_1t: in     vl_logic_vector(0 downto 0);
        seq_rdata_valid_lat_inc: out    vl_logic;
        seq_rdata_valid_lat_dec: out    vl_logic;
        ctl_rlat        : out    vl_logic_vector(4 downto 0);
        seq_poa_lat_dec_1x: out    vl_logic_vector(1 downto 0);
        seq_poa_lat_inc_1x: out    vl_logic_vector(1 downto 0);
        seq_poa_protection_override_1x: out    vl_logic;
        seq_oct_oct_delay: out    vl_logic_vector(4 downto 0);
        seq_oct_oct_extend: out    vl_logic_vector(4 downto 0);
        seq_oct_val     : out    vl_logic;
        seq_wdp_dqs_burst: out    vl_logic_vector(1 downto 0);
        seq_wdp_wdata_valid: out    vl_logic_vector(1 downto 0);
        seq_wdp_wdata   : out    vl_logic_vector(31 downto 0);
        seq_wdp_dm      : out    vl_logic_vector(3 downto 0);
        seq_wdp_dqs     : out    vl_logic_vector(1 downto 0);
        seq_wdp_ovride  : out    vl_logic;
        seq_dqs_add_2t_delay: out    vl_logic_vector(1 downto 0);
        ctl_wlat        : out    vl_logic_vector(4 downto 0);
        seq_mmc_start   : out    vl_logic;
        mmc_seq_done    : in     vl_logic;
        mmc_seq_value   : in     vl_logic;
        mem_err_out_n   : in     vl_logic;
        parity_error_n  : out    vl_logic;
        dbg_clk         : in     vl_logic;
        dbg_reset_n     : in     vl_logic;
        dbg_addr        : in     vl_logic_vector(12 downto 0);
        dbg_wr          : in     vl_logic;
        dbg_rd          : in     vl_logic;
        dbg_cs          : in     vl_logic;
        dbg_wr_data     : in     vl_logic_vector(31 downto 0);
        dbg_rd_data     : out    vl_logic_vector(31 downto 0);
        dbg_waitrequest : out    vl_logic
    );
end ddr2_phy_alt_mem_phy_seq_wrapper;
