library verilog;
use verilog.vl_types.all;
entity ddr2_phy_alt_mem_phy_addr_cmd is
    generic(
        DWIDTH_RATIO    : integer := 4;
        MEM_ADDR_CMD_BUS_COUNT: integer := 1;
        MEM_IF_BANKADDR_WIDTH: integer := 3;
        MEM_IF_CS_WIDTH : integer := 2;
        MEM_IF_MEMTYPE  : string  := "DDR";
        MEM_IF_ROWADDR_WIDTH: integer := 13
    );
    port(
        ac_clk_2x       : in     vl_logic;
        cs_n_clk_2x     : in     vl_logic;
        phy_clk_1x      : in     vl_logic;
        reset_ac_clk_2x_n: in     vl_logic;
        reset_cs_n_clk_2x_n: in     vl_logic;
        ctl_add_1t_ac_lat: in     vl_logic;
        ctl_add_1t_odt_lat: in     vl_logic;
        ctl_add_intermediate_regs: in     vl_logic;
        ctl_negedge_en  : in     vl_logic;
        ctl_mem_addr_h  : in     vl_logic_vector;
        ctl_mem_addr_l  : in     vl_logic_vector;
        ctl_mem_ba_h    : in     vl_logic_vector;
        ctl_mem_ba_l    : in     vl_logic_vector;
        ctl_mem_cas_n_h : in     vl_logic;
        ctl_mem_cas_n_l : in     vl_logic;
        ctl_mem_cke_h   : in     vl_logic_vector;
        ctl_mem_cke_l   : in     vl_logic_vector;
        ctl_mem_cs_n_h  : in     vl_logic_vector;
        ctl_mem_cs_n_l  : in     vl_logic_vector;
        ctl_mem_odt_h   : in     vl_logic_vector;
        ctl_mem_odt_l   : in     vl_logic_vector;
        ctl_mem_ras_n_h : in     vl_logic;
        ctl_mem_ras_n_l : in     vl_logic;
        ctl_mem_we_n_h  : in     vl_logic;
        ctl_mem_we_n_l  : in     vl_logic;
        seq_addr_h      : in     vl_logic_vector;
        seq_addr_l      : in     vl_logic_vector;
        seq_ba_h        : in     vl_logic_vector;
        seq_ba_l        : in     vl_logic_vector;
        seq_cas_n_h     : in     vl_logic;
        seq_cas_n_l     : in     vl_logic;
        seq_cke_h       : in     vl_logic_vector;
        seq_cke_l       : in     vl_logic_vector;
        seq_cs_n_h      : in     vl_logic_vector;
        seq_cs_n_l      : in     vl_logic_vector;
        seq_odt_h       : in     vl_logic_vector;
        seq_odt_l       : in     vl_logic_vector;
        seq_ras_n_h     : in     vl_logic;
        seq_ras_n_l     : in     vl_logic;
        seq_we_n_h      : in     vl_logic;
        seq_we_n_l      : in     vl_logic;
        seq_ac_sel      : in     vl_logic;
        mem_addr        : out    vl_logic_vector;
        mem_ba          : out    vl_logic_vector;
        mem_cas_n       : out    vl_logic;
        mem_cke         : out    vl_logic_vector;
        mem_cs_n        : out    vl_logic_vector;
        mem_odt         : out    vl_logic_vector;
        mem_ras_n       : out    vl_logic;
        mem_we_n        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADDR_CMD_BUS_COUNT : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_MEMTYPE : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ROWADDR_WIDTH : constant is 1;
end ddr2_phy_alt_mem_phy_addr_cmd;
