library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_input_if is
    generic(
        CFG_LOCAL_DATA_WIDTH: integer := 64;
        CFG_LOCAL_ID_WIDTH: integer := 8;
        CFG_LOCAL_ADDR_WIDTH: integer := 33;
        CFG_LOCAL_SIZE_WIDTH: integer := 3;
        CFG_MEM_IF_CHIP : integer := 1;
        CFG_AFI_INTF_PHASE_NUM: integer := 2;
        CFG_CTL_ARBITER_TYPE: string  := "ROWCOL"
    );
    port(
        itf_cmd_ready   : out    vl_logic;
        itf_cmd_valid   : in     vl_logic;
        itf_cmd         : in     vl_logic;
        itf_cmd_address : in     vl_logic_vector;
        itf_cmd_burstlen: in     vl_logic_vector;
        itf_cmd_id      : in     vl_logic_vector;
        itf_cmd_priority: in     vl_logic;
        itf_cmd_autopercharge: in     vl_logic;
        itf_cmd_multicast: in     vl_logic;
        itf_wr_data_ready: out    vl_logic;
        itf_wr_data_valid: in     vl_logic;
        itf_wr_data     : in     vl_logic_vector;
        itf_wr_data_byte_en: in     vl_logic_vector;
        itf_wr_data_begin: in     vl_logic;
        itf_wr_data_last: in     vl_logic;
        itf_wr_data_id  : in     vl_logic_vector;
        itf_rd_data_ready: in     vl_logic;
        itf_rd_data_valid: out    vl_logic;
        itf_rd_data     : out    vl_logic_vector;
        itf_rd_data_error: out    vl_logic;
        itf_rd_data_begin: out    vl_logic;
        itf_rd_data_last: out    vl_logic;
        itf_rd_data_id  : out    vl_logic_vector;
        itf_rd_data_id_early: out    vl_logic_vector;
        itf_rd_data_id_early_valid: out    vl_logic;
        cmd_gen_full    : in     vl_logic;
        cmd_valid       : out    vl_logic;
        cmd_address     : out    vl_logic_vector;
        cmd_write       : out    vl_logic;
        cmd_read        : out    vl_logic;
        cmd_multicast   : out    vl_logic;
        cmd_size        : out    vl_logic_vector;
        cmd_priority    : out    vl_logic;
        cmd_autoprecharge: out    vl_logic;
        cmd_id          : out    vl_logic_vector;
        wr_data_mem_full: in     vl_logic;
        write_data_id   : out    vl_logic_vector;
        write_data      : out    vl_logic_vector;
        byte_en         : out    vl_logic_vector;
        write_data_valid: out    vl_logic;
        read_data       : in     vl_logic_vector;
        read_data_valid : in     vl_logic;
        read_data_error : in     vl_logic;
        read_data_localid: in     vl_logic_vector;
        read_data_begin : in     vl_logic;
        read_data_last  : in     vl_logic;
        local_refresh_req: in     vl_logic;
        local_refresh_chip: in     vl_logic_vector;
        local_deep_powerdn_req: in     vl_logic;
        local_deep_powerdn_chip: in     vl_logic_vector;
        local_self_rfsh_req: in     vl_logic;
        local_self_rfsh_chip: in     vl_logic_vector;
        local_refresh_ack: out    vl_logic;
        local_deep_powerdn_ack: out    vl_logic;
        local_power_down_ack: out    vl_logic;
        local_self_rfsh_ack: out    vl_logic;
        local_init_done : out    vl_logic;
        bg_do_read      : in     vl_logic_vector;
        bg_do_rmw_correct: in     vl_logic_vector;
        bg_do_rmw_partial: in     vl_logic_vector;
        bg_localid      : in     vl_logic_vector;
        rfsh_req        : out    vl_logic;
        rfsh_chip       : out    vl_logic_vector;
        deep_powerdn_req: out    vl_logic;
        deep_powerdn_chip: out    vl_logic_vector;
        self_rfsh_req   : out    vl_logic;
        self_rfsh_chip  : out    vl_logic_vector;
        rfsh_ack        : in     vl_logic;
        deep_powerdn_ack: in     vl_logic;
        power_down_ack  : in     vl_logic;
        self_rfsh_ack   : in     vl_logic;
        init_done       : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_AFI_INTF_PHASE_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_CTL_ARBITER_TYPE : constant is 1;
end alt_mem_ddrx_input_if;
