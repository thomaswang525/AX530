`timescale 1ns / 1ps

module led_test (
                  clk,           // 开发板上输入时钟: 50Mhz
                  rst_n,         // 开发板上输入复位按键
                  led            // 输出LED灯,用于控制开发板上四个LED(LED1~LED4)
             );
             
//===========================================================================
// PORT declarations
//===========================================================================
input clk;
input rst_n;
output [3:0] led;

//寄存器定义
reg [31:0] timer;                  
reg [3:0] led;


//===========================================================================
// 计数器计数:循环计数0~4秒
//===========================================================================
  always @(posedge clk or negedge rst_n)    //检测时钟的上升沿和复位的下降沿
    begin
      if (~rst_n)                           //复位信号低有效
          timer <= 0;                       //计数器清零
      else if (timer == 32'd199_999_999)    //开发板使用的晶振为50MHz，4秒计数(50M*4-1=199_999_999)
          timer <= 0;                       //计数器计到4秒，计数器清零
      else
		    timer <= timer + 1'b1;            //计数器加1
    end

//===========================================================================
// LED灯控制
//===========================================================================
  always @(posedge clk or negedge rst_n)   //检测时钟的上升沿和复位的下降沿
    begin
      if (~rst_n)                          //复位信号低有效
          led <= 4'b1111;                  //LED灯输出全为高，四个LED灯灭           
      else if (timer == 32'd49_999_999)      //计数器计到1秒，
          led <= 4'b1110;                  //LED1点亮
      else if (timer == 32'd99_999_999)      //计数器计到2秒，
          led <= 4'b1101;                  //LED2点亮
      else if (timer == 32'd149_999_999)     //计数器计到3秒，
          led <= 4'b1011;                  //LED3点亮                           
      else if (timer == 32'd199_999_999)     //计数器计到4秒，
          led <= 4'b0111;                  //LED4点亮        
    end
    
endmodule

