library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_controller_st_top is
    generic(
        LOCAL_SIZE_WIDTH: string  := "";
        LOCAL_ADDR_WIDTH: string  := "";
        LOCAL_DATA_WIDTH: string  := "";
        LOCAL_BE_WIDTH  : string  := "";
        LOCAL_ID_WIDTH  : string  := "";
        LOCAL_CS_WIDTH  : string  := "";
        MEM_IF_ADDR_WIDTH: string  := "";
        MEM_IF_CLK_PAIR_COUNT: string  := "";
        LOCAL_IF_TYPE   : string  := "";
        DWIDTH_RATIO    : string  := "";
        CTL_ODT_ENABLED : string  := "";
        CTL_OUTPUT_REGD : string  := "";
        CTL_TBP_NUM     : string  := "";
        WRBUFFER_ADDR_WIDTH: string  := "";
        RDBUFFER_ADDR_WIDTH: string  := "";
        MEM_IF_CS_WIDTH : string  := "";
        MEM_IF_CHIP     : string  := "";
        MEM_IF_BANKADDR_WIDTH: string  := "";
        MEM_IF_ROW_WIDTH: string  := "";
        MEM_IF_COL_WIDTH: string  := "";
        MEM_IF_ODT_WIDTH: string  := "";
        MEM_IF_DQS_WIDTH: string  := "";
        MEM_IF_DWIDTH   : string  := "";
        MEM_IF_DM_WIDTH : string  := "";
        MAX_MEM_IF_CS_WIDTH: string  := "";
        MAX_MEM_IF_CHIP : string  := "";
        MAX_MEM_IF_BANKADDR_WIDTH: string  := "";
        MAX_MEM_IF_ROWADDR_WIDTH: string  := "";
        MAX_MEM_IF_COLADDR_WIDTH: string  := "";
        MAX_MEM_IF_ODT_WIDTH: string  := "";
        MAX_MEM_IF_DQS_WIDTH: string  := "";
        MAX_MEM_IF_DQ_WIDTH: string  := "";
        MAX_MEM_IF_MASK_WIDTH: string  := "";
        MAX_LOCAL_DATA_WIDTH: string  := "";
        CFG_TYPE        : string  := "";
        CFG_INTERFACE_WIDTH: string  := "";
        CFG_BURST_LENGTH: string  := "";
        CFG_DEVICE_WIDTH: string  := "";
        CFG_REORDER_DATA: string  := "";
        CFG_DATA_REORDERING_TYPE: string  := "";
        CFG_STARVE_LIMIT: string  := "";
        CFG_ADDR_ORDER  : string  := "";
        MEM_CAS_WR_LAT  : string  := "";
        MEM_ADD_LAT     : string  := "";
        MEM_TCL         : string  := "";
        MEM_TRRD        : string  := "";
        MEM_TFAW        : string  := "";
        MEM_TRFC        : string  := "";
        MEM_TREFI       : string  := "";
        MEM_TRCD        : string  := "";
        MEM_TRP         : string  := "";
        MEM_TWR         : string  := "";
        MEM_TWTR        : string  := "";
        MEM_TRTP        : string  := "";
        MEM_TRAS        : string  := "";
        MEM_TRC         : string  := "";
        CFG_TCCD        : string  := "";
        MEM_AUTO_PD_CYCLES: string  := "";
        CFG_SELF_RFSH_EXIT_CYCLES: string  := "";
        CFG_PDN_EXIT_CYCLES: string  := "";
        CFG_POWER_SAVING_EXIT_CYCLES: string  := "";
        CFG_MEM_CLK_ENTRY_CYCLES: string  := "";
        MEM_TMRD_CK     : string  := "";
        CTL_ECC_ENABLED : string  := "";
        CTL_ECC_RMW_ENABLED: string  := "";
        CTL_ECC_MULTIPLES_16_24_40_72: string  := "";
        CFG_GEN_SBE     : string  := "";
        CFG_GEN_DBE     : string  := "";
        CFG_ENABLE_INTR : string  := "";
        CFG_MASK_SBE_INTR: string  := "";
        CFG_MASK_DBE_INTR: string  := "";
        CFG_MASK_CORRDROP_INTR: integer := 0;
        CFG_CLR_INTR    : string  := "";
        CTL_USR_REFRESH : string  := "";
        CTL_REGDIMM_ENABLED: string  := "";
        CTL_ENABLE_BURST_INTERRUPT: string  := "";
        CTL_ENABLE_BURST_TERMINATE: string  := "";
        CFG_WRITE_ODT_CHIP: string  := "";
        CFG_READ_ODT_CHIP: string  := "";
        CFG_PORT_WIDTH_WRITE_ODT_CHIP: string  := "";
        CFG_PORT_WIDTH_READ_ODT_CHIP: string  := "";
        MEM_IF_CKE_WIDTH: string  := "";
        CTL_CSR_ENABLED : string  := "";
        CFG_ENABLE_NO_DM: string  := "";
        CSR_ADDR_WIDTH  : string  := "";
        CSR_DATA_WIDTH  : string  := "";
        CSR_BE_WIDTH    : string  := "";
        CFG_ENABLE_DQS_TRACKING: integer := 0;
        CFG_WLAT_BUS_WIDTH: integer := 6;
        CFG_RLAT_BUS_WIDTH: integer := 6;
        CFG_RRANK_BUS_WIDTH: integer := 0;
        CFG_WRANK_BUS_WIDTH: integer := 0;
        CFG_USE_SHADOW_REGS: integer := 0;
        MEM_IF_RD_TO_WR_TURNAROUND_OCT: string  := "";
        MEM_IF_WR_TO_RD_TURNAROUND_OCT: string  := "";
        CTL_RD_TO_PCH_EXTRA_CLK: integer := 0;
        CTL_RD_TO_RD_DIFF_CHIP_EXTRA_CLK: integer := 0;
        CTL_WR_TO_WR_DIFF_CHIP_EXTRA_CLK: integer := 0;
        CTL_ENABLE_WDATA_PATH_LATENCY: integer := 0;
        CFG_ECC_DECODER_REG: integer := 0;
        CFG_ERRCMD_FIFO_REG: integer := 0;
        ENABLE_BURST_MERGE: integer := 0
    );
    port(
        clk             : in     vl_logic;
        half_clk        : in     vl_logic;
        reset_n         : in     vl_logic;
        itf_cmd_ready   : out    vl_logic;
        itf_cmd_valid   : in     vl_logic;
        itf_cmd         : in     vl_logic;
        itf_cmd_address : in     vl_logic_vector;
        itf_cmd_burstlen: in     vl_logic_vector;
        itf_cmd_id      : in     vl_logic_vector;
        itf_cmd_priority: in     vl_logic;
        itf_cmd_autopercharge: in     vl_logic;
        itf_cmd_multicast: in     vl_logic;
        itf_wr_data_ready: out    vl_logic;
        itf_wr_data_valid: in     vl_logic;
        itf_wr_data     : in     vl_logic_vector;
        itf_wr_data_byte_en: in     vl_logic_vector;
        itf_wr_data_begin: in     vl_logic;
        itf_wr_data_last: in     vl_logic;
        itf_wr_data_id  : in     vl_logic_vector;
        itf_rd_data_ready: in     vl_logic;
        itf_rd_data_valid: out    vl_logic;
        itf_rd_data     : out    vl_logic_vector;
        itf_rd_data_error: out    vl_logic;
        itf_rd_data_begin: out    vl_logic;
        itf_rd_data_last: out    vl_logic;
        itf_rd_data_id  : out    vl_logic_vector;
        afi_rst_n       : out    vl_logic_vector;
        afi_cs_n        : out    vl_logic_vector;
        afi_cke         : out    vl_logic_vector;
        afi_odt         : out    vl_logic_vector;
        afi_addr        : out    vl_logic_vector;
        afi_ba          : out    vl_logic_vector;
        afi_ras_n       : out    vl_logic_vector;
        afi_cas_n       : out    vl_logic_vector;
        afi_we_n        : out    vl_logic_vector;
        afi_dqs_burst   : out    vl_logic_vector;
        afi_wdata_valid : out    vl_logic_vector;
        afi_wdata       : out    vl_logic_vector;
        afi_dm          : out    vl_logic_vector;
        afi_wlat        : in     vl_logic_vector;
        afi_rdata_en    : out    vl_logic_vector;
        afi_rdata_en_full: out    vl_logic_vector;
        afi_rdata       : in     vl_logic_vector;
        afi_rdata_valid : in     vl_logic_vector;
        afi_rrank       : out    vl_logic_vector;
        afi_wrank       : out    vl_logic_vector;
        afi_rlat        : in     vl_logic_vector;
        afi_cal_success : in     vl_logic;
        afi_cal_fail    : in     vl_logic;
        afi_cal_req     : out    vl_logic;
        afi_init_req    : out    vl_logic;
        afi_mem_clk_disable: out    vl_logic_vector;
        afi_cal_byte_lane_sel_n: out    vl_logic_vector;
        afi_ctl_refresh_done: out    vl_logic_vector;
        afi_seq_busy    : in     vl_logic_vector;
        afi_ctl_long_idle: out    vl_logic_vector;
        local_init_done : out    vl_logic;
        local_refresh_ack: out    vl_logic;
        local_powerdn_ack: out    vl_logic;
        local_self_rfsh_ack: out    vl_logic;
        local_deep_powerdn_ack: out    vl_logic;
        local_refresh_req: in     vl_logic;
        local_refresh_chip: in     vl_logic_vector;
        local_powerdn_req: in     vl_logic;
        local_self_rfsh_req: in     vl_logic;
        local_self_rfsh_chip: in     vl_logic_vector;
        local_deep_powerdn_req: in     vl_logic;
        local_deep_powerdn_chip: in     vl_logic_vector;
        local_multicast : in     vl_logic;
        local_priority  : in     vl_logic;
        ecc_interrupt   : out    vl_logic;
        csr_read_req    : in     vl_logic;
        csr_write_req   : in     vl_logic;
        csr_burst_count : in     vl_logic_vector(0 downto 0);
        csr_beginbursttransfer: in     vl_logic;
        csr_addr        : in     vl_logic_vector;
        csr_wdata       : in     vl_logic_vector;
        csr_rdata       : out    vl_logic_vector;
        csr_be          : in     vl_logic_vector;
        csr_rdata_valid : out    vl_logic;
        csr_waitrequest : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOCAL_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_BE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CLK_PAIR_COUNT : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_IF_TYPE : constant is 1;
    attribute mti_svvh_generic_type of DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CTL_ODT_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_OUTPUT_REGD : constant is 1;
    attribute mti_svvh_generic_type of CTL_TBP_NUM : constant is 1;
    attribute mti_svvh_generic_type of WRBUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of RDBUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_ROWADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_COLADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_MASK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_INTERFACE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_BURST_LENGTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DEVICE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_REORDER_DATA : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_REORDERING_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_STARVE_LIMIT : constant is 1;
    attribute mti_svvh_generic_type of CFG_ADDR_ORDER : constant is 1;
    attribute mti_svvh_generic_type of MEM_CAS_WR_LAT : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADD_LAT : constant is 1;
    attribute mti_svvh_generic_type of MEM_TCL : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRRD : constant is 1;
    attribute mti_svvh_generic_type of MEM_TFAW : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRFC : constant is 1;
    attribute mti_svvh_generic_type of MEM_TREFI : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRCD : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRP : constant is 1;
    attribute mti_svvh_generic_type of MEM_TWR : constant is 1;
    attribute mti_svvh_generic_type of MEM_TWTR : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRTP : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRAS : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRC : constant is 1;
    attribute mti_svvh_generic_type of CFG_TCCD : constant is 1;
    attribute mti_svvh_generic_type of MEM_AUTO_PD_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_SELF_RFSH_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PDN_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_POWER_SAVING_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_CLK_ENTRY_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of MEM_TMRD_CK : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_RMW_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_MULTIPLES_16_24_40_72 : constant is 1;
    attribute mti_svvh_generic_type of CFG_GEN_SBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_GEN_DBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_MASK_SBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_MASK_DBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_MASK_CORRDROP_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_CLR_INTR : constant is 1;
    attribute mti_svvh_generic_type of CTL_USR_REFRESH : constant is 1;
    attribute mti_svvh_generic_type of CTL_REGDIMM_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_ENABLE_BURST_INTERRUPT : constant is 1;
    attribute mti_svvh_generic_type of CTL_ENABLE_BURST_TERMINATE : constant is 1;
    attribute mti_svvh_generic_type of CFG_WRITE_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_READ_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_WRITE_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_READ_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CKE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CTL_CSR_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_NO_DM : constant is 1;
    attribute mti_svvh_generic_type of CSR_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CSR_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CSR_BE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_DQS_TRACKING : constant is 1;
    attribute mti_svvh_generic_type of CFG_WLAT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_RLAT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_RRANK_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_WRANK_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_USE_SHADOW_REGS : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_RD_TO_WR_TURNAROUND_OCT : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_WR_TO_RD_TURNAROUND_OCT : constant is 1;
    attribute mti_svvh_generic_type of CTL_RD_TO_PCH_EXTRA_CLK : constant is 1;
    attribute mti_svvh_generic_type of CTL_RD_TO_RD_DIFF_CHIP_EXTRA_CLK : constant is 1;
    attribute mti_svvh_generic_type of CTL_WR_TO_WR_DIFF_CHIP_EXTRA_CLK : constant is 1;
    attribute mti_svvh_generic_type of CTL_ENABLE_WDATA_PATH_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_DECODER_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ERRCMD_FIFO_REG : constant is 1;
    attribute mti_svvh_generic_type of ENABLE_BURST_MERGE : constant is 1;
end alt_mem_ddrx_controller_st_top;
