library verilog;
use verilog.vl_types.all;
entity ddr2_alt_mem_ddrx_controller_top is
    port(
        clk             : in     vl_logic;
        half_clk        : in     vl_logic;
        reset_n         : in     vl_logic;
        local_ready     : out    vl_logic;
        local_write     : in     vl_logic;
        local_read      : in     vl_logic;
        local_address   : in     vl_logic_vector(24 downto 0);
        local_byteenable: in     vl_logic_vector(3 downto 0);
        local_writedata : in     vl_logic_vector(31 downto 0);
        local_burstcount: in     vl_logic_vector(2 downto 0);
        local_beginbursttransfer: in     vl_logic;
        local_readdata  : out    vl_logic_vector(31 downto 0);
        local_readdatavalid: out    vl_logic;
        afi_rst_n       : out    vl_logic_vector(0 downto 0);
        afi_cs_n        : out    vl_logic_vector(0 downto 0);
        afi_cke         : out    vl_logic_vector(0 downto 0);
        afi_odt         : out    vl_logic_vector(0 downto 0);
        afi_addr        : out    vl_logic_vector(12 downto 0);
        afi_ba          : out    vl_logic_vector(2 downto 0);
        afi_ras_n       : out    vl_logic_vector(0 downto 0);
        afi_cas_n       : out    vl_logic_vector(0 downto 0);
        afi_we_n        : out    vl_logic_vector(0 downto 0);
        afi_dqs_burst   : out    vl_logic_vector(1 downto 0);
        afi_wdata_valid : out    vl_logic_vector(1 downto 0);
        afi_wdata       : out    vl_logic_vector(31 downto 0);
        afi_dm          : out    vl_logic_vector(3 downto 0);
        afi_wlat        : in     vl_logic_vector(4 downto 0);
        afi_rdata_en    : out    vl_logic_vector(1 downto 0);
        afi_rdata_en_full: out    vl_logic_vector(1 downto 0);
        afi_rdata       : in     vl_logic_vector(31 downto 0);
        afi_rdata_valid : in     vl_logic_vector(0 downto 0);
        afi_rlat        : in     vl_logic_vector(4 downto 0);
        afi_cal_success : in     vl_logic;
        afi_cal_fail    : in     vl_logic;
        afi_cal_req     : out    vl_logic;
        afi_mem_clk_disable: out    vl_logic_vector(0 downto 0);
        afi_cal_byte_lane_sel_n: out    vl_logic_vector(1 downto 0);
        afi_ctl_refresh_done: out    vl_logic_vector(0 downto 0);
        afi_seq_busy    : in     vl_logic_vector(0 downto 0);
        afi_ctl_long_idle: out    vl_logic_vector(0 downto 0);
        local_init_done : out    vl_logic;
        local_refresh_ack: out    vl_logic;
        local_powerdn_ack: out    vl_logic;
        local_self_rfsh_ack: out    vl_logic;
        local_autopch_req: in     vl_logic;
        local_refresh_req: in     vl_logic;
        local_refresh_chip: in     vl_logic_vector(0 downto 0);
        local_powerdn_req: in     vl_logic;
        local_self_rfsh_req: in     vl_logic;
        local_self_rfsh_chip: in     vl_logic_vector(0 downto 0);
        local_multicast : in     vl_logic;
        local_priority  : in     vl_logic;
        ecc_interrupt   : out    vl_logic;
        csr_read_req    : in     vl_logic;
        csr_write_req   : in     vl_logic;
        csr_burst_count : in     vl_logic_vector(0 downto 0);
        csr_beginbursttransfer: in     vl_logic;
        csr_addr        : in     vl_logic_vector(15 downto 0);
        csr_wdata       : in     vl_logic_vector(31 downto 0);
        csr_rdata       : out    vl_logic_vector(31 downto 0);
        csr_be          : in     vl_logic_vector(3 downto 0);
        csr_rdata_valid : out    vl_logic;
        csr_waitrequest : out    vl_logic
    );
end ddr2_alt_mem_ddrx_controller_top;
